module task1(input [9:0]sw, output [9:0]led);
	assign led = sw;
endmodule
